module writeback_mux #(
    parameter W = 32
)(
    input logic [W-1:0] ReadData,
    input logic [W-1:0] ALUResult,
    input logic ResultSrc,

    output logic [W-1:0] Result
)