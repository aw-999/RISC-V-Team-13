module ControlUnit #(
    parameter AD = 5
)(
    input logic [6:0] opcode,
    input logic [14:12] funct3,
    input logic funct7,

    //flags
    input logic Zero,
    input logic Negative,

    output logic RegWriteD,
    output logic
    output logic
    output logic
    output logic
    output logic
    output logic
    output logic
    


)